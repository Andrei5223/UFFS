library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entidade principal
ENTITY BN IS
    PORT(
        escolha_jogador : IN STD_LOGIC_VECTOR(3 downto 0);  -- Escolha do jogador
        codificacao_barco_inserido : IN STD_LOGIC_VECTOR(4 downto 0); -- Codifica��o do barco sendo inserido
        barco: IN STD_LOGIC_VECTOR(2 downto 0); --Escolhe qual barco est� inserindo
        clock: IN STD_LOGIC
    );
END BN;


-- Cria tabuleiro
ARCHITECTURE Behavior_Tabuleiro OF BN IS 

                                    -- �ndices da matriz (3 em inteiro)            -- Conte�do do �ndice (vetor de 4 bits)
    TYPE matriz_tabuleiro IS ARRAY (natural range 0 to 3, natural range 0 to 3) of std_logic_vector(3 downto 0);
    SIGNAL matriz : matriz_tabuleiro;   -- Cria matriz

BEGIN

    --Salvar a 
    PROCESS (clock)

    --Para salvar a codifica��o das posi��es escolhidas
	variable pos1 : STD_LOGIC_VECTOR(3 downto 0);
	variable pos2: STD_LOGIC_VECTOR(3 downto 0);
	variable pos3 : STD_LOGIC_VECTOR(3 downto 0);
	variable pos4: STD_LOGIC_VECTOR(3 downto 0);

    BEGIN
    matriz(0, 0) <= "0110";
    matriz(0, 1) <= "1101";
    matriz(0, 2) <= "1000";
    matriz(0, 3) <= "0011";
    matriz(1, 0) <= "0000";
    matriz(1, 1) <= "1001";
    matriz(1, 2) <= "0001";
    matriz(1, 3) <= "1011";
    matriz(2, 0) <= "0111";
    matriz(2, 1) <= "0100";
    matriz(2, 2) <= "1110";
    matriz(2, 3) <= "0010";
    matriz(3, 0) <= "0101";
    matriz(3, 1) <= "1111";
    matriz(3, 2) <= "1010";
    matriz(3, 3) <= "1100";

    END PROCESS;
END Behavior_Tabuleiro;